library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity control_memory_20332993 is
    Port ( IN_CAR : in std_logic_vector(16 downto 0);
           FL : out std_logic; -- 0
           RZ : out std_logic; -- 1
           RN : out std_logic; -- 2
           RC : out std_logic; -- 3
           RV : out std_logic; -- 4
           MW : out std_logic; -- 5
           MM : out std_logic; -- 6
           RW : out std_logic; -- 7
           MD : out std_logic; -- 8
           FS : out std_logic_vector(4 downto 0); -- 9 to 13
           MB : out std_logic; -- 14
           TB : out std_logic; -- 15
           TA : out std_logic; -- 16
           TD : out std_logic; -- 17
           PL : out std_logic; -- 18
           PI : out std_logic; -- 19
           IL : out std_logic; -- 20
           MC : out std_logic; -- 21
           MS : out std_logic_vector(2 downto 0); -- 22 to 24
           NA : out std_logic_vector(16 downto 0) -- 25 to 41
    );
end control_memory_20332993;

architecture Behavioral of control_memory_20332993 is

-- we will use the least significant 8 bit of the IN_CAR - array(0 to 255)
type mem_array is array(0 to 255) of std_logic_vector(41 downto 0);
-- initialise the control memory
signal control_mem : mem_array := (
 -- |41 25|2422|21|20|19|18|17|16|15|14|13 9|8|7|6|5|4|3|2|1|0|
 -- | Next Address | MS | M| I| P| P| T| T| T| M| FS |M|R|M|M|R|R|R|R|F|
 -- | Next Address | MS | C| L| I| L| D| A| B| B| FS |D|W|M|W|V|C|N|Z|L|
 -- "00000000000000000 000 0 0 0 0 0 0 0 0 00000 0 0 0 0 0 0 0 0 0"

    "000000000010111010000000000000000111000000", --Load values into first 32 registers
    "000000000010111100000000100000000111000000", --Load value into the 33rd register
  --"000000000000000000000000100000000111000000"
 --                              |||||
    "000000000010111110000000000000100010000000", --A + not B
    "000000000011000000000000000001010010000000", --A or B
    "000000000011000010000000000000011010000000", --A + B + 1
    "000000000011000100000000000001100010000000", --A xor B
    "000000000011000110000000000000010010000000", --A + B 
    "000000000011001000000000000011000010000000", --sl B
    "000000000011001010000000000000000010000000", --A 
    "000000000011001100000000000010000010000000", --B
    "000000000011001110000000000000001010000000", --A + 1
    "000000000011010000000000000000101010000000", --A + not B + 1
    "000000000011010010000000000000110010000000", --A - 1
    "000000000011010100000000000001110010000000", --not A
    "000000000011010110000000000001000010000000", --A & B
    "000000000011011000000000000010100010000000", --sr B
    "000000000011011010000000000000111010000000", --A
    "000000000011011100000000000000000000000000", 
    "000000000011011110000000000000000000000000", 
    "000000000011100000000000000000000000000000",
    "000000000011100010000000000000000000000000",
    "000000000011100100000000000000000000000000",
    "000000000011100110000000000000000000000000",
    "000000000011101000000000000000000000000000", "000000000011101010000000000000000000000000", "000000000011101100000000000000000000000000", "000000000011101110000000000000000000000000", "000000000011110000000000000000000000000000", "000000000011110010000000000000000000000000", "000000000011110100000000000000000000000000", "000000000011110110000000000000000000000000", "000000000011111000000000000000000000000000", "000000000011111010000000000000000000000000", "000000000011111100000000000000000000000000", "000000000011111110000000000000000000000000", "000000000100000000000000000000000000000000", "000000000100000010000000000000000000000000", "000000000100000100000000000000000000000000", "000000000100000110000000000000000000000000", "000000000100001000000000000000000000000000", "000000000100001010000000000000000000000000", "000000000100001100000000000000000000000000", "000000000100001110000000000000000000000000", "000000000100010000000000000000000000000000", "000000000100010010000000000000000000000000", "000000000100010100000000000000000000000000", "000000000100010110000000000000000000000000", "000000000100011000000000000000000000000000", "000000000100011010000000000000000000000000", "000000000100011100000000000000000000000000", "000000000100011110000000000000000000000000", "000000000100100000000000000000000000000000", "000000000100100010000000000000000000000000", "000000000100100100000000000000000000000000", "000000000100100110000000000000000000000000", "000000000100101000000000000000000000000000", "000000000100101010000000000000000000000000", "000000000100101100000000000000000000000000", "000000000100101110000000000000000000000000", "000000000100110000000000000000000000000000", "000000000100110010000000000000000000000000", "000000000100110100000000000000000000000000", "000000000100110110000000000000000000000000", "000000000100111000000000000000000000000000", "000000000100111010000000000000000000000000", "000000000100111100000000000000000000000000", "000000000100111110000000000000000000000000", "000000000101000000000000000000000000000000", "000000000101000010000000000000000000000000", "000000000101000100000000000000000000000000", "000000000101000110000000000000000000000000", "000000000101001000000000000000000000000000", "000000000101001010000000000000000000000000", "000000000101001100000000000000000000000000", "000000000101001110000000000000000000000000", "000000000101010000000000000000000000000000", "000000000101010010000000000000000000000000", "000000000101010100000000000000000000000000", "000000000101010110000000000000000000000000", "000000000101011000000000000000000000000000", "000000000101011010000000000000000000000000", "000000000101011100000000000000000000000000", "000000000101011110000000000000000000000000", "000000000101100000000000000000000000000000", "000000000101100010000000000000000000000000", "000000000101100100000000000000000000000000", "000000000101100110000000000000000000000000", "000000000101101000000000000000000000000000", "000000000101101010000000000000000000000000", "000000000101101100000000000000000000000000", "000000000101101110000000000000000000000000", "000000000101110000000000000000000000000000", "000000000101110010000000000000000000000000", "000000000101110100000000000000000000000000", "000000000101110110000000000000000000000000", "000000000101111000000000000000000000000000", "000000000101111010000000000000000000000000", "000000000101111100000000000000000000000000", "000000000101111110000000000000000000000000", "000000000110000000000000000000000000000000", "000000000110000010000000000000000000000000", "000000000110000100000000000000000000000000", "000000000110000110000000000000000000000000", "000000000110001000000000000000000000000000", "000000000110001010000000000000000000000000", "000000000110001100000000000000000000000000", "000000000110001110000000000000000000000000", "000000000110010000000000000000000000000000", "000000000110010010000000000000000000000000", "000000000110010100000000000000000000000000", "000000000110010110000000000000000000000000", "000000000110011000000000000000000000000000", "000000000110011010000000000000000000000000", "000000000110011100000000000000000000000000", "000000000110011110000000000000000000000000", "000000000110100000000000000000000000000000", "000000000110100010000000000000000000000000", "000000000110100100000000000000000000000000", "000000000110100110000000000000000000000000", "000000000110101000000000000000000000000000", "000000000110101010000000000000000000000000", "000000000110101100000000000000000000000000", "000000000110101110000000000000000000000000", "000000000110110000000000000000000000000000", "000000000110110010000000000000000000000000", "000000000110110100000000000000000000000000", "000000000110110110000000000000000000000000", "000000000110111000000000000000000000000000", "000000000110111010000000000000000000000000", "000000000110111100000000000000000000000000", "000000000110111110000000000000000000000000", "000000000111000000000000000000000000000000", "000000000111000010000000000000000000000000", "000000000111000100000000000000000000000000", "000000000111000110000000000000000000000000", "000000000111001000000000000000000000000000", "000000000111001010000000000000000000000000", "000000000111001100000000000000000000000000", "000000000111001110000000000000000000000000", "000000000111010000000000000000000000000000", "000000000111010010000000000000000000000000", "000000000111010100000000000000000000000000", "000000000111010110000000000000000000000000", "000000000111011000000000000000000000000000", "000000000111011010000000000000000000000000", "000000000111011100000000000000000000000000", "000000000111011110000000000000000000000000", "000000000111100000000000000000000000000000", "000000000111100010000000000000000000000000", "000000000111100100000000000000000000000000", "000000000111100110000000000000000000000000", "000000000111101000000000000000000000000000", "000000000111101010000000000000000000000000", "000000000111101100000000000000000000000000", "000000000111101110000000000000000000000000", "000000000111110000000000000000000000000000", "000000000111110010000000000000000000000000", "000000000111110100000000000000000000000000", "000000000111110110000000000000000000000000", "000000000111111000000000000000000000000000", "000000000111111010000000000000000000000000", "000000000111111100000000000000000000000000", "000000000111111110000000000000000000000000", "000000001000000000000000000000000000000000", "000000001000000010000000000000000000000000", "000000001000000100000000000000000000000000", "000000001000000110000000000000000000000000", "000000001000001000000000000000000000000000", "000000001000001010000000000000000000000000", "000000001000001100000000000000000000000000", "000000001000001110000000000000000000000000", "000000001000010000000000000000000000000000", "000000001000010010000000000000000000000000", "000000001000010100000000000000000000000000", "000000001000010110000000000000000000000000", "000000001000011000000000000000000000000000", "000000001000011010000000000000000000000000", "000000001000011100000000000000000000000000", "000000001000011110000000000000000000000000", "000000001000100000000000000000000000000000", "000000001000100010000000000000000000000000", "000000001000100100000000000000000000000000", "000000001000100110000000000000000000000000", "000000001000101000000000000000000000000000", "000000001000101010000000000000000000000000", "000000001000101100000000000000000000000000", "000000001000101110000000000000000000000000", "000000001000110000000000000000000000000000", "000000001000110010000000000000000000000000", "000000001000110100000000000000000000000000", "000000001000110110000000000000000000000000", "000000001000111000000000000000000000000000", "000000001000111010000000000000000000000000", "000000001000111100000000000000000000000000", "000000001000111110000000000000000000000000", "000000001001000000000000000000000000000000", "000000001001000010000000000000000000000000", "000000001001000100000000000000000000000000", "000000001001000110000000000000000000000000", "000000001001001000000000000000000000000000", "000000001001001010000000000000000000000000", "000000001001001100000000000000000000000000", "000000001001001110000000000000000000000000", "000000001001010000000000000000000000000000", "000000001001010010000000000000000000000000", "000000001001010100000000000000000000000000", "000000001001010110000000000000000000000000", "000000001001011000000000000000000000000000", "000000001001011010000000000000000000000000", "000000001001011100000000000000000000000000", "000000001001011110000000000000000000000000", "000000001001100000000000000000000000000000", "000000001001100010000000000000000000000000", "000000001001100100000000000000000000000000", "000000001001100110000000000000000000000000", "000000001001101000000000000000000000000000", "000000001001101010000000000000000000000000", "000000001001101100000000000000000000000000", "000000001001101110000000000000000000000000", "000000001001110000000000000000000000000000", "000000001001110010000000000000000000000000", "000000001001110100000000000000000000000000", "000000001001110110000000000000000000000000", "000000001001111000000000000000000000000000", "000000001001111010000000000000000000000000", "000000001001111100000000000000000000000000", "000000001001111110000000000000000000000000", "000000001010000000000000000000000000000000", "000000001010000010000000000000000000000000", "000000001010000100000000000000000000000000", "000000001010000110000000000000000000000000", "000000001010001000000000000000000000000000", "000000001010001010000000000000000000000000", "000000001010001100000000000000000000000000", "000000001010001110000000000000000000000000", "000000001010010000000000000000000000000000", "000000001010010010000000000000000000000000", "000000001010010100000000000000000000000000", "000000001010010110000000000000000000000000", "000000001010011000000000000000000000000000", "000000001010011010000000000000000000000000", "000000001010011100000000000000000000000000", "000000001010011110000000000000000000000000", "000000001010100000000000000000000000000000", "000000001010100010000000000000000000000000", "000000001010100100000000000000000000000000", "000000001010100110000000000000000000000000", "000000001010101000000000000000000000000000", "000000001010101010000000000000000000000000", "000000001010101100000000000000000000000000", "000000001010101110000000000000000000000000", "000000001010110000000000000000000000000000", "000000001010110010000000000000000000000000", "000000001010110100000000000000000000000000", "000000001010110110000000000000000000000000", "000000001010111000000000000000000000000000" 
);

signal content_at_address : std_logic_vector(41 downto 0); 

begin
    content_at_address <= control_mem(to_integer(unsigned(IN_CAR(8 downto 0)))) after 2ns;
    FL <= content_at_address(0); -- 0
    RZ <= content_at_address(1); -- 1
    RN <= content_at_address(2); -- 2
    RC <= content_at_address(3); -- 3
    RV <= content_at_address(4); -- 4
    MW <= content_at_address(5); -- 5
    MM <= content_at_address(6); -- 6
    RW <= content_at_address(7); -- 7
    MD <= content_at_address(8); -- 8
    FS <= content_at_address(13 downto 9); -- 9 to 13
    MB <= content_at_address(14); -- 14
    TB <= content_at_address(15); -- 15
    TA <= content_at_address(16); -- 16
    TD <= content_at_address(17); -- 17
    PL <= content_at_address(18); -- 18
    PI <= content_at_address(19); -- 19
    IL <= content_at_address(20); -- 20
    MC <= content_at_address(21); -- 21
    MS <= content_at_address(24 downto 22); -- 22 to 24
    NA <= content_at_address(41 downto 25); -- 25 to 41

end Behavioral;
