library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity memory_module_20332993 is
  Port (address : in std_logic_vector(31 downto 0);
        write_data : in std_logic_vector(31 downto 0);
        write_enable : in std_logic;
        clock : in std_logic;
        read_data : out std_logic_vector(31 downto 0));
end memory_module_20332993;

architecture Behavioral of memory_module_20332993 is
  -- we will use the least significant 4 bit of the address - array(0 to 16)
  type mem_array is array(0 to 511) of std_logic_vector(31 downto 0);
  -- initialize data memory, X denotes hexadecimal numberend Behavioral;
  signal data_mem : mem_array := (
  X"00000000", X"00000001", X"00000002", X"00000003", X"00000004", X"00000005", X"00000006", X"00000007", X"00000008", X"00000009", X"0000000a", X"0000000b", X"0000000c", X"0000000d", X"0000000e", X"0000000f", X"00000010", X"00000011", X"00000012", X"00000013", X"00000014", X"00000015", X"00000016", X"00000017", X"00000018", X"00000019", X"0000001a", X"0000001b", X"0000001c", X"0000001d", X"0000001e", X"0000001f", X"00000020", X"00000021", X"00000022", X"00000023", X"00000024", X"00000025", X"00000026", X"00000027", X"00000028", X"00000029", X"0000002a", X"0000002b", X"0000002c", X"0000002d", X"0000002e", X"0000002f", X"00000030", X"00000031", X"00000032", X"00000033", X"00000034", X"00000035", X"00000036", X"00000037", X"00000038", X"00000039", X"0000003a", X"0000003b", X"0000003c", X"0000003d", X"0000003e", X"0000003f", X"00000040", X"00000041", X"00000042", X"00000043", X"00000044", X"00000045", X"00000046", X"00000047", X"00000048", X"00000049", X"0000004a", X"0000004b", X"0000004c", X"0000004d", X"0000004e", X"0000004f", X"00000050", X"00000051", X"00000052", X"00000053", X"00000054", X"00000055", X"00000056", X"00000057", X"00000058", X"00000059", X"0000005a", X"0000005b", X"0000005c", X"0000005d", X"0000005e", X"0000005f", X"00000060", X"00000061", X"00000062", X"00000063", X"00000064", X"00000065", X"00000066", X"00000067", X"00000068", X"00000069", X"0000006a", X"0000006b", X"0000006c", X"0000006d", X"0000006e", X"0000006f", X"00000070", X"00000071", X"00000072", X"00000073", X"00000074", X"00000075", X"00000076", X"00000077", X"00000078", X"00000079", X"0000007a", X"0000007b", X"0000007c", X"0000007d", X"0000007e", X"0000007f", X"00000080", X"00000081", X"00000082", X"00000083", X"00000084", X"00000085", X"00000086", X"00000087", X"00000088", X"00000089", X"0000008a", X"0000008b", X"0000008c", X"0000008d", X"0000008e", X"0000008f", X"00000090", X"00000091", X"00000092", X"00000093", X"00000094", X"00000095", X"00000096", X"00000097", X"00000098", X"00000099", X"0000009a", X"0000009b", X"0000009c", X"0000009d", X"0000009e", X"0000009f", X"000000a0", X"000000a1", X"000000a2", X"000000a3", X"000000a4", X"000000a5", X"000000a6", X"000000a7", X"000000a8", X"000000a9", X"000000aa", X"000000ab", X"000000ac", X"000000ad", X"000000ae", X"000000af", X"000000b0", X"000000b1", X"000000b2", X"000000b3", X"000000b4", X"000000b5", X"000000b6", X"000000b7", X"000000b8", X"000000b9", X"000000ba", X"000000bb", X"000000bc", X"000000bd", X"000000be", X"000000bf", X"000000c0", X"000000c1", X"000000c2", X"000000c3", X"000000c4", X"000000c5", X"000000c6", X"000000c7", X"000000c8", X"000000c9", X"000000ca", X"000000cb", X"000000cc", X"000000cd", X"000000ce", X"000000cf", X"000000d0", X"000000d1", X"000000d2", X"000000d3", X"000000d4", X"000000d5", X"000000d6", X"000000d7", X"000000d8", X"000000d9", X"000000da", X"000000db", X"000000dc", X"000000dd", X"000000de", X"000000df", X"000000e0", X"000000e1", X"000000e2", X"000000e3", X"000000e4", X"000000e5", X"000000e6", X"000000e7", X"000000e8", X"000000e9", X"000000ea", X"000000eb", X"000000ec", X"000000ed", X"000000ee", X"000000ef", X"000000f0", X"000000f1", X"000000f2", X"000000f3", X"000000f4", X"000000f5", X"000000f6", X"000000f7", X"000000f8", X"000000f9", X"000000fa", X"000000fb", X"000000fc", X"000000fd", X"000000fe", X"000000ff", X"00000100", X"00000101", X"00000102", X"00000103", X"00000104", X"00000105", X"00000106", X"00000107", X"00000108", X"00000109", X"0000010a", X"0000010b", X"0000010c", X"0000010d", X"0000010e", X"0000010f", X"00000110", X"00000111", X"00000112", X"00000113", X"00000114", X"00000115", X"00000116", X"00000117", X"00000118", X"00000119", X"0000011a", X"0000011b", X"0000011c", X"0000011d", X"0000011e", X"0000011f", X"00000120", X"00000121", X"00000122", X"00000123", X"00000124", X"00000125", X"00000126", X"00000127", X"00000128", X"00000129", X"0000012a", X"0000012b", X"0000012c", X"0000012d", X"0000012e", X"0000012f", X"00000130", X"00000131", X"00000132", X"00000133", X"00000134", X"00000135", X"00000136", X"00000137", X"00000138", X"00000139", X"0000013a", X"0000013b", X"0000013c", X"0000013d", X"0000013e", X"0000013f", X"00000140", X"00000141", X"00000142", X"00000143", X"00000144", X"00000145", X"00000146", X"00000147", X"00000148", X"00000149", X"0000014a", X"0000014b", X"0000014c", X"0000014d", X"0000014e", X"0000014f", X"00000150", X"00000151", X"00000152", X"00000153", X"00000154", X"00000155", X"00000156", X"00000157", X"00000158", X"00000159", X"0000015a", X"0000015b", X"0000015c", X"0000015d", X"0000015e", X"0000015f", X"00000160", X"00000161", X"00000162", X"00000163", X"00000164", X"00000165", X"00000166", X"00000167", X"00000168", X"00000169", X"0000016a", X"0000016b", X"0000016c", X"0000016d", X"0000016e", X"0000016f", X"00000170", X"00000171", X"00000172", X"00000173", X"00000174", X"00000175", X"00000176", X"00000177", X"00000178", X"00000179", X"0000017a", X"0000017b", X"0000017c", X"0000017d", X"0000017e", X"0000017f", X"00000180", X"00000181", X"00000182", X"00000183", X"00000184", X"00000185", X"00000186", X"00000187", X"00000188", X"00000189", X"0000018a", X"0000018b", X"0000018c", X"0000018d", X"0000018e", X"0000018f", X"00000190", X"00000191", X"00000192", X"00000193", X"00000194", X"00000195", X"00000196", X"00000197", X"00000198", X"00000199", X"0000019a", X"0000019b", X"0000019c", X"0000019d", X"0000019e", X"0000019f", X"000001a0", X"000001a1", X"000001a2", X"000001a3", X"000001a4", X"000001a5", X"000001a6", X"000001a7", X"000001a8", X"000001a9", X"000001aa", X"000001ab", X"000001ac", X"000001ad", X"000001ae", X"000001af", X"000001b0", X"000001b1", X"000001b2", X"000001b3", X"000001b4", X"000001b5", X"000001b6", X"000001b7", X"000001b8", X"000001b9", X"000001ba", X"000001bb", X"000001bc", X"000001bd", X"000001be", X"000001bf", X"000001c0", X"000001c1", X"000001c2", X"000001c3", X"000001c4", X"000001c5", X"000001c6", X"000001c7", X"000001c8", X"000001c9", X"000001ca", X"000001cb", X"000001cc", X"000001cd", X"000001ce", X"000001cf", X"000001d0", X"000001d1", X"000001d2", X"000001d3", X"000001d4", X"000001d5", X"000001d6", X"000001d7", X"000001d8", X"000001d9", X"000001da", X"000001db", X"000001dc", X"000001dd", X"000001de", X"000001df", X"000001e0", X"000001e1", X"000001e2", X"000001e3", X"000001e4", X"000001e5", X"000001e6", X"000001e7", X"000001e8", X"000001e9", X"000001ea", X"000001eb", X"000001ec", X"000001ed", X"000001ee", X"000001ef", X"000001f0", X"000001f1", X"000001f2", X"000001f3", X"000001f4", X"000001f5", X"000001f6", X"000001f7", X"000001f8", X"000001f9", X"000001fa", X"000001fb", X"000001fc", X"000001fd", X"000001fe", X"000001ff"
  );
begin
mem_process: process(clock)
begin
  if(rising_edge(clock)) then
    if(write_enable='1') then
      data_mem(to_integer(unsigned(address(8 downto 0)))) <= write_data after 2ns;
    end if;
  end if;
end process;
read_data <= data_mem(to_integer(unsigned(address(8 downto 0)))) after 2ns;
end Behavioral;
