library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity decoder_6to32_20332993 is
    Port (  S : in  std_logic_vector (4 downto 0);
            Extra : in std_logic;
            z : out std_logic_vector(31 downto 0));
end decoder_6to32_20332993;

architecture Behavioral of decoder_6to32_20332993 is

begin

process (S, Extra)
    begin
    if(Extra='1') then
      z <= "00000000000000000000000000000000";
    else     
    case S is
      when "00000" => z <= "00000000000000000000000000000001"; 
      when "00001" => z <= "00000000000000000000000000000010";
      when "00010" => z <= "00000000000000000000000000000100";
      when "00011" => z <= "00000000000000000000000000001000";
      when "00100" => z <= "00000000000000000000000000010000";
      when "00101" => z <= "00000000000000000000000000100000";
      when "00110" => z <= "00000000000000000000000001000000";
      when "00111" => z <= "00000000000000000000000010000000";
      when "01000" => z <= "00000000000000000000000100000000";
      when "01001" => z <= "00000000000000000000001000000000";
      when "01010" => z <= "00000000000000000000010000000000";
      when "01011" => z <= "00000000000000000000100000000000";
      when "01100" => z <= "00000000000000000001000000000000";
      when "01101" => z <= "00000000000000000010000000000000";
      when "01110" => z <= "00000000000000000100000000000000";
      when "01111" => z <= "00000000000000001000000000000000";
      when "10000" => z <= "00000000000000010000000000000000";
      when "10001" => z <= "00000000000000100000000000000000";
      when "10010" => z <= "00000000000001000000000000000000";
      when "10011" => z <= "00000000000010000000000000000000";
      when "10100" => z <= "00000000000100000000000000000000";
      when "10101" => z <= "00000000001000000000000000000000";
      when "10110" => z <= "00000000010000000000000000000000";
      when "10111" => z <= "00000000100000000000000000000000";
      when "11000" => z <= "00000001000000000000000000000000";
      when "11001" => z <= "00000010000000000000000000000000";
      when "11010" => z <= "00000100000000000000000000000000";
      when "11011" => z <= "00001000000000000000000000000000";
      when "11100" => z <= "00010000000000000000000000000000";
      when "11101" => z <= "00100000000000000000000000000000";
      when "11110" => z <= "01000000000000000000000000000000";
      when "11111" => z <= "10000000000000000000000000000000";
      when others => z <= "00000000000000000000000000000000";
    end case;
    end if;
  end process;

end Behavioral;
